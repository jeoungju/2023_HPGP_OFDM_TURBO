`timescale 1ps/1ps
module testbench();

parameter D_WIDTH = 4;
parameter A_WIDTH = 9;
parameter COS_SIN = 16;


reg clk, n_rst;
reg start;
reg mode_3072_384;
reg in_vld;
reg [3:0] in_re, in_im;

wire [6:0] out_re, out_im;
wire out_vld;


always #5 clk = ~clk;
    initial begin
        clk = 1'b0;
        n_rst = 1'b0;
        #7 n_rst = 1'b1;
    end

initial begin
    start = 1'b0;
    mode_3072_384 = 1'b0;
    in_vld = 1'b0;
    in_re = 4'h0;
    in_im = 4'h0;
    #33;
    start = 1'b1;
    mode_3072_384 = 1'b1;
    in_vld = 1'b1;
    in_re = 4'h1;
    in_im = 4'h0;
    #90;
    in_re = 4'h4;
    in_im = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'h4;
    #10;




    $stop;
end

/*
initial begin
    start = 1'b0;
    mode_3072_384 = 1'b0;
    in_vld = 1'b0;
    in_re = 4'h0;
    in_im = 4'h0;
    #33;
    start = 1'b1;
    mode_3072_384 = 1'b1;
    in_vld = 1'b1;
    in_re = 4'h1;
    in_im = 4'h0;
    #90;
    in_re = 4'h4;
    in_im = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;
    in_re = 4'hc;
    #10;
    in_re = 4'h4;
    #10;



    $stop;
end
*/
full_384 dut_full_384(
    .clk(clk),
	.n_rst(n_rst),
	.start(start),
    .mode_3072_384(mode_3072_384),
	.in_vld(in_vld),
	.in_re(in_re),
	.in_im(in_re),
	.out_re(out_re),
	.out_im(out_im),
	.out_vld(out_vld)
);

endmodule
