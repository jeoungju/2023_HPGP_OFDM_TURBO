`timescale 1ns/100ps
`define T_CLK 10
module testbench;

reg clk, n_rst;


parameter D1_SIZE = 13;
parameter D2_SIZE = 11;
parameter SIGN_BIT=1;
parameter INT_BIT=6;
parameter FLT_BIT=6;


reg [D1_SIZE-1:0] in1_re, in1_im;
reg [D1_SIZE-1:0] in2_re, in2_im;
reg [D1_SIZE-1:0] in3_re, in3_im;

wire [D1_SIZE+1:0] out1_re, out1_im;
wire [D1_SIZE+1:0] out2_re, out2_im;
wire [D1_SIZE+1:0] out3_re, out3_im;

reg din_vld;
wire dout_vld;



always #5 clk = ~clk;
    initial begin
        clk = 1'b0;
        n_rst = 1'b0;
        #7 n_rst = 1'b1;
    end

/////////BOUNDARY CONDITION ////////////
// 13'b1_000_010_000_000; //-62
// 13'b0_111_110_000_000; // 62
// 13'b0_100_001_000_000; // 33
// 13'b0_011_111_000_000; // 31
// 13'b0_000_001_000_000; //  1
// 13'b0_000_010_000_000; //  2
// 13'b1_111_110_000_000; // -2
// 13'b1_111_111_000_000; // -1
/////////////////////////////////////////

initial begin
	din_vld = 1'b0;
	in1_re = 0;
	in1_im = 0;
	in2_re = 0;
	in2_im = 0;
	in3_re = 0;
	in3_im = 0;

	#33;

//case1_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b0_000_001_000_000; //1
	in1_im = 13'b0_000_001_000_000; //1
	in2_re = 13'b0_000_010_000_000; //2
	in2_im = 13'b0_000_010_000_000; //2
	in3_re = 13'b1_111_111_000_000; //-1
	in3_im = 13'b1_111_111_000_000; //-1
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case1_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b0_000_001_000_000; //1
	in2_im = 13'b0_000_001_000_000; //1
	in1_re = 13'b0_000_010_000_000; //2
	in1_im = 13'b0_000_010_000_000; //2
	in3_re = 13'b1_111_111_000_000; //-1
	in3_im = 13'b1_111_111_000_000; //-1
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case2_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b1_000_010_000_000; //-62
	in1_im = 13'b1_000_010_000_000; //-62
	in2_re = 13'b0_000_010_000_000; //2
	in2_im = 13'b0_000_010_000_000; //2
	in3_re = 13'b0_011_111_000_000;// 31
	in3_im = 13'b0_011_111_000_000; // 31
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case2_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b1_000_010_000_000; //-62
	in2_im = 13'b1_000_010_000_000; //-62
	in1_re = 13'b0_000_010_000_000; //2
	in1_im = 13'b0_000_010_000_000; //2
	in3_re = 13'b0_011_111_000_000; // 31
	in3_im = 13'b0_011_111_000_000; // 31
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case2_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b1_000_010_000_000; //-62
	in3_im = 13'b1_000_010_000_000; //-62
	in2_re = 13'b0_000_010_000_000; //2
	in2_im = 13'b0_000_010_000_000; //2
	in1_re = 13'b0_011_111_000_000; // 31
	in1_im = 13'b0_011_111_000_000; // 31
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case3_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b0_011_111_000_000; // 31
	in1_im = 13'b0_011_111_000_000; // 31
	in2_re = 13'b0_100_001_000_000; // 33
	in2_im = 13'b0_100_001_000_000; // 33
	in3_re = 13'b0_111_110_000_000; // 62
	in3_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case3_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b0_011_111_000_000; // 31
	in2_im = 13'b0_011_111_000_000; // 31
	in1_re = 13'b0_100_001_000_000; // 33
	in1_im = 13'b0_100_001_000_000; // 33
	in3_re = 13'b0_111_110_000_000; // 62
	in3_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case3_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b0_011_111_000_000; // 31
	in3_im = 13'b0_011_111_000_000; // 31
	in2_re = 13'b0_100_001_000_000; // 33
	in2_im = 13'b0_100_001_000_000; // 33
	in1_re = 13'b0_111_110_000_000; // 62
	in1_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case4_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b1_111_110_000_000; // -2
	in1_im = 13'b1_111_110_000_000; // -2
	in2_re = 13'b1_000_010_000_000; //-62
	in2_im = 13'b1_000_010_000_000; //-62
	in3_re = 13'b0_111_110_000_000; // 62
	in3_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case4_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b1_111_110_000_000; // -2
	in2_im = 13'b1_111_110_000_000; // -2
	in1_re = 13'b1_000_010_000_000; //-62
	in1_im = 13'b1_000_010_000_000;//-62
	in3_re = 13'b0_111_110_000_000;// 62
	in3_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case4_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b1_111_110_000_000; // -2
	in3_im = 13'b1_111_110_000_000; // -2
	in2_re = 13'b1_000_010_000_000; //-62
	in2_im = 13'b1_000_010_000_000; //-62
	in1_re = 13'b0_111_110_000_000; // 62
	in1_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case5_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b0_011_111_000_000; // 31
	in1_im = 13'b0_011_111_000_000; // 31
	in2_re = 13'b0_100_001_000_000; // 33
	in2_im = 13'b0_100_001_000_000; // 33
	in3_re = 13'b0_111_110_000_000; // 62
	in3_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case5_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b0_011_111_000_000; // 31
	in2_im = 13'b0_011_111_000_000; // 31
	in1_re = 13'b0_100_001_000_000; // 33
	in1_im = 13'b0_100_001_000_000; // 33
	in3_re = 13'b0_111_110_000_000;// 62
	in3_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case5_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b0_011_111_000_000; // 31
	in3_im = 13'b0_011_111_000_000; // 31
	in2_re = 13'b0_100_001_000_000; // 33
	in2_im = 13'b0_100_001_000_000; // 33
	in1_re = 13'b0_111_110_000_000; // 62
	in1_im = 13'b0_111_110_000_000; // 62
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case6_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b1_111_110_000_000; //-2
	in1_im = 13'b1_111_110_000_000; //-2
	in2_re = 13'b1_111_111_000_000; //-1
	in2_im = 13'b1_111_111_000_000; //-1
	in3_re = 13'b0_011_111_000_000; //31
	in3_im = 13'b0_011_111_000_000; //31
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case6_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b1_111_110_000_000; //-2
	in2_im = 13'b1_111_110_000_000; //-2
	in1_re = 13'b1_111_111_000_000; //-1
	in1_im = 13'b1_111_111_000_000; //-1
	in3_re = 13'b0_011_111_000_000; //31
	in3_im = 13'b0_011_111_000_000; //31
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case6_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b1_111_110_000_000; //-2
	in3_im = 13'b1_111_110_000_000; //-2
	in2_re = 13'b1_111_111_000_000; //-1
	in2_im = 13'b1_111_111_000_000; //-1
	in1_re = 13'b0_011_111_000_000; //31
	in1_im = 13'b0_011_111_000_000; //31
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case7_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b0_011_111_000_000; //31
	in1_im = 13'b0_011_111_000_000; //31
	in2_re = 13'b0_000_010_000_000; //2
	in2_im = 13'b0_000_010_000_000; //2
	in3_re = 13'b0_000_001_000_000; //1
	in3_im = 13'b0_000_001_000_000; //1
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case7_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b0_011_111_000_000; //31
	in2_im = 13'b0_011_111_000_000; //31
	in1_re = 13'b0_000_010_000_000; //2
	in1_im = 13'b0_000_010_000_000; //2
	in3_re = 13'b0_000_001_000_000; //1
	in3_im = 13'b0_000_001_000_000; //1
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case7_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b0_011_111_000_000; //31
	in3_im = 13'b0_011_111_000_000; //31
	in2_re = 13'b0_000_010_000_000; //2
	in2_im = 13'b0_000_010_000_000; //2
	in1_re = 13'b0_000_001_000_000; //1
	in1_im = 13'b0_000_001_000_000; //1
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case8_1
/////////////////////////////////////////
	din_vld = 1'b1;
	in1_re = 13'b0_000_010_000_000; //2
	in1_im = 13'b0_000_010_000_000; //2
	in2_re = 13'b1_111_110_000_000; //-2
	in2_im = 13'b1_111_110_000_000; //-2
	in3_re = 13'b0_000_010_000_000; //2
	in3_im = 13'b0_000_010_000_000; //2
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case8_2
/////////////////////////////////////////
	din_vld = 1'b1;
	in2_re = 13'b0_000_010_000_000; //2
	in2_im = 13'b0_000_010_000_000; //2
	in1_re = 13'b1_111_110_000_000; //-2
	in1_im = 13'b1_111_110_000_000; //-2
	in3_re = 13'b0_000_010_000_000; //2
	in3_im = 13'b0_000_010_000_000; //2
	#10;
	din_vld = 1'b0;
	#50;
/////////////////////////////////////////
//case8_3
/////////////////////////////////////////
	din_vld = 1'b1;
	in3_re = 13'b0_000_010_000_000; //2
	in3_im = 13'b0_000_010_000_000; //2
	in2_re = 13'b1_111_110_000_000; //-2
	in2_im = 13'b1_111_110_000_000; //-2
	in1_re = 13'b0_000_010_000_000; //2
	in1_im = 13'b0_000_010_000_000; //2
	#10;
	din_vld = 1'b0;
	#100;
/////////////////////////////////////////
//case9_1
/////////////////////////////////////////
din_vld = 1'b1;
in1_re = 13'b0_111_110_000_000; //62
in1_im = 13'b0_111_110_000_000; //62
in2_re = 13'b1_000_010_000_000; //-62
in2_im = 13'b1_000_010_000_000; //-62
in3_re = 13'b0_000_101_000_000; //5
in3_im = 13'b0_000_101_000_000; //5
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case9_2
/////////////////////////////////////////
din_vld = 1'b1;
in2_re = 13'b0_111_110_000_000; //62
in2_im = 13'b0_111_110_000_000; //62
in1_re = 13'b1_000_010_000_000; //-62
in1_im = 13'b1_000_010_000_000; //-62
in3_re = 13'b0_000_101_000_000; //5
in3_im = 13'b0_000_101_000_000; //5
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case9_3
/////////////////////////////////////////
din_vld = 1'b1;
in3_re = 13'b0_111_110_000_000; //62
in3_im = 13'b0_111_110_000_000; //62
in2_re = 13'b1_000_010_000_000; //-62
in2_im = 13'b1_000_010_000_000; //-62
in1_re = 13'b0_000_101_000_000; //5
in1_im = 13'b0_000_101_000_000; //5
#10;
din_vld = 1'b0;
#100;
/////////////////////////////////////////
//case10_1
/////////////////////////////////////////
din_vld = 1'b1;
in1_re = 13'b0_000_111_000_000; //7
in1_im = 13'b0_000_111_000_000; //7
in2_re = 13'b0_100_001_000_000; // 33
in2_im = 13'b0_100_001_000_000; // 33
in3_re = 13'b1_111_111_000_000; //-1
in3_im = 13'b1_111_111_000_000; //-1
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case10_2
/////////////////////////////////////////
din_vld = 1'b1;
in2_re = 13'b0_000_111_000_000; //7
in2_im = 13'b0_000_111_000_000; //7
in1_re = 13'b0_100_001_000_000; // 33
in1_im = 13'b0_100_001_000_000; // 33
in3_re = 13'b1_111_111_000_000; //-1
in3_im = 13'b1_111_111_000_000; //-1
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case10_3
/////////////////////////////////////////
din_vld = 1'b1;
in3_re = 13'b0_000_111_000_000; //7
in3_im = 13'b0_000_111_000_000; //7
in2_re = 13'b0_100_001_000_000; // 33
in2_im = 13'b0_100_001_000_000; // 33
in1_re = 13'b1_111_111_000_000; //-1
in1_im = 13'b1_111_111_000_000; //-1
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case11_1
/////////////////////////////////////////
din_vld = 1'b1;
in1_re = 13'b0_100_001_000_000; // 33
in1_im = 13'b0_100_001_000_000; // 33
in2_re = 13'b0_001_010_000_000; //10
in2_im = 13'b0_001_010_000_000; //10
in3_re = 13'b0_111_110_000_000; //62
in3_im = 13'b0_111_110_000_000; //62
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case11_2
/////////////////////////////////////////
din_vld = 1'b1;
in2_re = 13'b0_100_001_000_000; // 33
in2_im = 13'b0_100_001_000_000; // 33
in1_re = 13'b0_001_010_000_000; //10
in1_im = 13'b0_001_010_000_000; //10
in3_re = 13'b0_111_110_000_000; //62
in3_im = 13'b0_111_110_000_000; //62
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////
//case11_3
/////////////////////////////////////////
din_vld = 1'b1;
in3_re = 13'b0_100_001_000_000; // 33
in3_im = 13'b0_100_001_000_000; // 33
in2_re = 13'b0_001_010_000_000; //10
in2_im = 13'b0_001_010_000_000; //10
in1_re = 13'b0_111_110_000_000; //62
in1_im = 13'b0_111_110_000_000; //62
#10;
din_vld = 1'b0;
#50;
/////////////////////////////////////////


	$stop;

end

rd3bf #(
    .SIGN_BIT(SIGN_BIT),
    .INT_BIT(INT_BIT),
    .FLT_BIT(FLT_BIT)
) u_rd3bf (
	.clk(clk),
	.n_rst(n_rst),
	.di_vld(din_vld),
	.in1_re(in1_re), 
	.in1_im(in1_im),
    .in2_re(in2_re), 
	.in2_im(in2_im),
    .in3_re(in3_re), 
	.in3_im(in3_im),
	.out1_re(out1_re), 
	.out1_im(out1_im),
    .out2_re(out2_re), 
	.out2_im(out2_im),
    .out3_re(out3_re), 
	.out3_im(out3_im),
	.do_vld(dout_vld)
);


endmodule
